`timescale 1ns / 1ps

// Complete program testbench for Vigna RISC-V processor
// Tests complete C programs compiled to RISC-V machine code

module program_testbench();

    // Clock and reset
    reg clk;
    reg resetn;
    
    // Instruction memory interface
    wire        i_valid;
    reg         i_ready;
    wire [31:0] i_addr;
    reg  [31:0] i_rdata;
    
    // Data memory interface  
    wire        d_valid;
    reg         d_ready;
    wire [31:0] d_addr;
    reg  [31:0] d_rdata;
    wire [31:0] d_wdata;
    wire [ 3:0] d_wstrb;
    
    // Test control
    reg [31:0] instruction_memory [0:1023];
    reg [31:0] data_memory [0:1023];
    integer test_pass_count;
    integer test_fail_count;
    integer cycle_count;
    reg [31:0] last_pc;
    integer same_pc_count;
    
    // Expected test results for verification
    integer expected_fib[8];
    integer expected_sorted[5];
    
    // Instantiate the processor core
    vigna dut (
        .clk(clk),
        .resetn(resetn),
        .i_valid(i_valid),
        .i_ready(i_ready),
        .i_addr(i_addr),
        .i_rdata(i_rdata),
        .d_valid(d_valid),
        .d_ready(d_ready),
        .d_addr(d_addr),
        .d_rdata(d_rdata),
        .d_wdata(d_wdata),
        .d_wstrb(d_wstrb)
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    // Instruction memory simulation
    always @(posedge clk) begin
        if (resetn) begin
            if (i_valid && !i_ready) begin
                i_rdata <= instruction_memory[i_addr[11:2]];
                i_ready <= 1;
            end else begin
                i_ready <= 0;
            end
        end else begin
            i_ready <= 0;
        end
    end
    
    // Data memory simulation
    always @(posedge clk) begin
        if (resetn) begin
            if (d_valid && !d_ready) begin
                if (d_wstrb != 0) begin
                    // Write operation
                    // Map address 0x1000+ to data_memory starting at index 0
                    if (d_wstrb == 4'b1111) begin
                        data_memory[(d_addr - 32'h1000) >> 2] <= d_wdata;
                        // $display("DEBUG: Write to addr=0x%08x, data=0x%08x, mem_idx=%d", d_addr, d_wdata, (d_addr - 32'h1000) >> 2);
                    end else if (d_wstrb == 4'b0011)
                        data_memory[(d_addr - 32'h1000) >> 2] <= (data_memory[(d_addr - 32'h1000) >> 2] & 32'hFFFF0000) | (d_wdata & 32'h0000FFFF);
                    else if (d_wstrb == 4'b0001)
                        data_memory[(d_addr - 32'h1000) >> 2] <= (data_memory[(d_addr - 32'h1000) >> 2] & 32'hFFFFFF00) | (d_wdata & 32'h000000FF);
                end else begin
                    // Read operation
                    d_rdata <= data_memory[(d_addr - 32'h1000) >> 2];
                end
                d_ready <= 1;
            end else begin
                d_ready <= 0;
            end
        end else begin
            d_ready <= 0;
        end
    end
    
    // Load specific program into instruction memory
    task load_simple_test;
        begin
            $display("Loading simple_test program...");
            // Clear memory
            for (integer i = 0; i < 1024; i = i + 1) begin
                instruction_memory[i] = 32'h00000013; // NOP
                data_memory[i] = 32'h00000000;
            end
            
            // Load program - include the generated assignments
            `include "programs/build/simple_test.vh"
            $display("Simple test program loaded successfully");
        end
    endtask
    
    task load_fibonacci_test;
        begin
            $display("Loading fibonacci_simple program...");
            // Clear memory
            for (integer i = 0; i < 1024; i = i + 1) begin
                instruction_memory[i] = 32'h00000013; // NOP
                data_memory[i] = 32'h00000000;
            end
            
            // Load program - include the generated assignments
            `include "programs/build/fibonacci_simple.vh"
            $display("Fibonacci simple program loaded successfully");
        end
    endtask
    
    // Run program with timeout
    task run_program;
        input [255:0] test_name;
        input integer max_cycles;
        
        begin
            $display("Running program: %s", test_name);
            
            cycle_count = 0;
            last_pc = 32'hFFFFFFFF;
            same_pc_count = 0;
            
            while (cycle_count < max_cycles) begin
                @(posedge clk);
                cycle_count = cycle_count + 1;
                
                // Check for infinite loop (same PC for multiple cycles)
                if (i_addr == last_pc) begin
                    same_pc_count = same_pc_count + 1;
                    if (same_pc_count >= 10) begin
                        $display("Program halted at PC=0x%08x after %d cycles", i_addr, cycle_count);
                        cycle_count = max_cycles; // Exit loop
                    end
                end else begin
                    same_pc_count = 0;
                    last_pc = i_addr;
                end
            end
            
            if (same_pc_count < 10) begin
                $display("Program timeout after %d cycles", max_cycles);
            end
        end
    endtask
    
    // Verify test results
    task verify_simple_test_results;
        integer base_addr;
        begin
            $display("Verifying simple test results...");
            
            // Check result at data_memory[0x1000/4] = data_memory[1024]
            // But our data memory is only 1024 words, so check at base of our range
            // The program writes to 0x1000, 0x1004, 0x1008, 0x100C
            // We'll check data_memory[0x1000>>2] which is outside our range
            // Let's adjust the test to write to lower addresses by modifying our expectation
            
            $display("Data memory contents:");
            for (integer i = 0; i < 8; i = i + 1) begin
                if (data_memory[i] != 0) begin
                    $display("  data_memory[%d] = 0x%08x (%d)", i, data_memory[i], data_memory[i]);
                end
            end
            
            // The program writes to addresses 0x1000, 0x1004, 0x1008, 0x100C
            // With our address mapping, these map to data_memory[0], [1], [2], [3]
            base_addr = 0;
            
            if (base_addr < 1024) begin
                // Check first result: should be 30 (10 + 20)
                if (data_memory[base_addr] == 32'd30) begin
                    $display("  PASS: Arithmetic test result = %d (expected 30)", data_memory[base_addr]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: Arithmetic test result = %d (expected 30)", data_memory[base_addr]);
                    test_fail_count = test_fail_count + 1;
                end
                
                // Check second result: should be 15 (1+2+3+4+5)
                if (data_memory[base_addr + 1] == 32'd15) begin
                    $display("  PASS: Loop test result = %d (expected 15)", data_memory[base_addr + 1]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: Loop test result = %d (expected 15)", data_memory[base_addr + 1]);
                    test_fail_count = test_fail_count + 1;
                end
                
                // Check third result: should be 20 (max of 10, 20)
                if (data_memory[base_addr + 2] == 32'd20) begin
                    $display("  PASS: Conditional test result = %d (expected 20)", data_memory[base_addr + 2]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: Conditional test result = %d (expected 20)", data_memory[base_addr + 2]);
                    test_fail_count = test_fail_count + 1;
                end
                
                // Check completion marker: should be 0xDEADBEEF
                if (data_memory[base_addr + 3] == 32'hDEADBEEF) begin
                    $display("  PASS: Completion marker = 0x%08x (expected 0xDEADBEEF)", data_memory[base_addr + 3]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: Completion marker = 0x%08x (expected 0xDEADBEEF)", data_memory[base_addr + 3]);
                    test_fail_count = test_fail_count + 1;
                end
            end else begin
                $display("  FAIL: Program writes to addresses outside our data memory range");
                test_fail_count = test_fail_count + 4;
            end
        end
    endtask
    
    // Verify fibonacci test results
    task verify_fibonacci_test_results;
        integer base_addr;
        begin
            $display("Verifying fibonacci test results...");
            base_addr = 0;
            
            // Expected Fibonacci sequence: 0, 1, 1, 2, 3, 5, 8, 13
            
            for (integer i = 0; i < 8; i = i + 1) begin
                if (data_memory[base_addr + i] == expected_fib[i]) begin
                    $display("  PASS: fib[%d] = %d (expected %d)", i, data_memory[base_addr + i], expected_fib[i]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: fib[%d] = %d (expected %d)", i, data_memory[base_addr + i], expected_fib[i]);
                    test_fail_count = test_fail_count + 1;
                end
            end
            
            // Check completion marker
            if (data_memory[base_addr + 8] == 32'h12345678) begin
                $display("  PASS: Completion marker = 0x%08x (expected 0x12345678)", data_memory[base_addr + 8]);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: Completion marker = 0x%08x (expected 0x12345678)", data_memory[base_addr + 8]);
                test_fail_count = test_fail_count + 1;
            end
        end
    endtask
    
    // Verify sorting test results
    task verify_sorting_test_results;
        integer base_addr;
        begin
            $display("Verifying sorting test results...");
            base_addr = 0;
            
            // Expected sorted array: {1, 2, 5, 8, 9} (from original {5, 2, 8, 1, 9})
            
            for (integer i = 0; i < 5; i = i + 1) begin
                if (data_memory[base_addr + i] == expected_sorted[i]) begin
                    $display("  PASS: sorted[%d] = %d (expected %d)", i, data_memory[base_addr + i], expected_sorted[i]);
                    test_pass_count = test_pass_count + 1;
                end else begin
                    $display("  FAIL: sorted[%d] = %d (expected %d)", i, data_memory[base_addr + i], expected_sorted[i]);
                    test_fail_count = test_fail_count + 1;
                end
            end
            
            // Check completion marker
            if (data_memory[base_addr + 5] == 32'hABCDEF00) begin
                $display("  PASS: Completion marker = 0x%08x (expected 0xABCDEF00)", data_memory[base_addr + 5]);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: Completion marker = 0x%08x (expected 0xABCDEF00)", data_memory[base_addr + 5]);
                test_fail_count = test_fail_count + 1;
            end
        end
    endtask
    
    // Main test sequence
    initial begin
        $dumpfile("program_test.vcd");
        $dumpvars(0, program_testbench);
        
        $display("Starting Complete Program Tests for Vigna Processor");
        $display("=================================================");
        
        // Initialize
        resetn = 0;
        test_pass_count = 0;
        test_fail_count = 0;
        
        // Initialize expected results
        expected_fib[0] = 0;
        expected_fib[1] = 1;
        expected_fib[2] = 1;
        expected_fib[3] = 2;
        expected_fib[4] = 3;
        expected_fib[5] = 5;
        expected_fib[6] = 8;
        expected_fib[7] = 13;
        
        expected_sorted[0] = 1;
        expected_sorted[1] = 2;
        expected_sorted[2] = 5;
        expected_sorted[3] = 8;
        expected_sorted[4] = 9;
        
        // Reset pulse
        repeat(10) @(posedge clk);
        resetn = 1;
        
        // Test 1: Simple arithmetic program
        load_simple_test();
        run_program("Simple Arithmetic Test", 1000);
        verify_simple_test_results();
        
        // Reset processor between tests
        $display("");
        $display("Resetting processor for next test...");
        resetn = 0;
        repeat(10) @(posedge clk);
        resetn = 1;
        
        // Test 2: Fibonacci program
        $display("");
        load_fibonacci_test();
        run_program("Fibonacci Test", 3000);
        verify_fibonacci_test_results();
        
        // Test summary
        $display("");
        $display("Complete Program Test Summary:");
        $display("=============================");
        $display("Tests Passed: %d", test_pass_count);
        $display("Tests Failed: %d", test_fail_count);
        $display("Total Tests:  %d", test_pass_count + test_fail_count);
        
        if (test_fail_count == 0) begin
            $display("All complete program tests PASSED!");
        end else begin
            $display("Some complete program tests FAILED!");
        end
        
        $finish;
    end

endmodule