//////////////////////////////////////////////////////////////////////////////////
// Company: Wuhan University
// Engineer: Xuanyu Hu
// 
// Create Date: 2022/04/27 16:39:33
// Design Name: vigna_v1
// Module Name: vigna
// Project Name: vigna
// Description: A simple RV32I CPU core
// 
// Dependencies: none
// 
// Revision: 
// Revision 1.09
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifndef VIGNA_CORE_V 
`define VIGNA_CORE_V

`timescale 1ns / 1ps
`include "vigna_conf.vh"

`ifdef VIGNA_CORE_M_EXTENSION
`include "vigna_coproc.v"
`endif 

//vigna top module
module vigna(
    input clk,
    input resetn,

`ifdef VIGNA_CORE_INTERRUPT
    // Interrupt inputs
    input             ext_irq,      // External interrupt
    input             timer_irq,    // Timer interrupt
    input             soft_irq,     // Software interrupt
`endif

    output            i_valid,
    input             i_ready,
    output     [31:0] i_addr,
    input      [31:0] i_rdata,

    output reg        d_valid,
    input             d_ready,
    output reg [31:0] d_addr,
    input      [31:0] d_rdata,
    output reg [31:0] d_wdata,
    output reg [ 3:0] d_wstrb
);

//program counter
reg  [31:0] pc;
wire [31:0] pc_next;

//part 1: fetching unit
reg  [31:0] inst;
wire [31:0] inst_addr;
reg  [ 1:0] fetch_state;
reg  internal_valid;

`ifdef VIGNA_CORE_C_EXTENSION
reg  [15:0] pending_inst; // Store upper 16 bits when fetching compressed instruction
reg  inst_is_16bit;       // Flag indicating current instruction is 16-bit
reg  have_pending;        // Flag indicating we have a pending upper 16 bits  
`endif

wire fetched, fetch_received;
assign fetched = fetch_state == 3;



//assign inst = i_ready ? i_rdata : inst;
assign inst_addr = i_addr;
assign i_addr = pc;

assign i_valid = internal_valid;

always @ (posedge clk) begin
    //reset logic
    if (!resetn) begin
        pc              <= `VIGNA_CORE_RESET_ADDR;
        fetch_state     <= 0;
        internal_valid  <= 0;
        `ifdef VIGNA_CORE_C_EXTENSION
        pending_inst    <= 16'h0;
        inst_is_16bit   <= 0;
        have_pending    <= 0;
        `endif
    end else begin
        //fetch logic
        case (fetch_state)
            0: begin
                internal_valid     <= 1;
                fetch_state <= 1;
            end
            1: begin
                if (i_ready) begin
                    `ifdef VIGNA_CORE_C_EXTENSION
                    // Simple approach: check if lower 16 bits are compressed
                    if (i_rdata[1:0] != 2'b11) begin
                        // 16-bit compressed instruction
                        inst[31:16]   <= 16'h0;
                        inst[15:0]    <= i_rdata[15:0];
                        inst_is_16bit <= 1;
                    end else begin
                        // 32-bit instruction
                        inst          <= i_rdata;
                        inst_is_16bit <= 0;
                    end
                    `else
                    inst            <= i_rdata;
                    `endif
                    internal_valid  <= 0;
                    fetch_state     <= 3;
                end
            end
            3: begin
                if (fetch_received) begin
                    internal_valid  <= 1;
                    pc              <= pc_next;
                    fetch_state     <= 1;
                end
            end
            default: begin
                internal_valid  <= 0;
                fetch_state     <= 0;
            end
        endcase
    end
end

//decode logic
wire [6:0] opcode;
wire [2:0] funct3;
wire [6:0] funct7;
wire [4:0] rd;
wire [4:0] rs1;
wire [4:0] rs2;

assign opcode = effective_inst[6:0];
assign funct3 = effective_inst[14:12];
assign funct7 = effective_inst[31:25];
assign rd     = effective_inst[11:7];
assign rs1    = effective_inst[19:15];
assign rs2    = effective_inst[24:20];

//r
wire is_add, is_sub, is_sll, is_slt, is_sltu, is_xor, is_srl, is_sra, is_or, is_and;
//i
wire is_addi, is_slli, is_slti, is_sltiu, is_xori, is_srli, is_srai, is_ori, is_andi;
wire is_jalr, is_lb, is_lh, is_lw, is_lbu, is_lhu;
//s
wire is_sb, is_sh, is_sw;
//b
wire is_beq, is_bne, is_blt, is_bge, is_bltu, is_bgeu;
//u
wire is_lui, is_auipc;
//j
wire is_jal;

wire funct7_zero, funct7_sub_sra;
assign funct7_zero = funct7 == 0;
assign funct7_sub_sra = funct7 == 7'b0100000;

wire i_type_alu, i_type_jalr, i_type_load;
assign i_type_alu  = opcode == 7'b0010011;
assign i_type_jalr = opcode == 7'b1100111;
assign i_type_load = opcode == 7'b0000011;

`ifdef VIGNA_CORE_ZICSR_EXTENSION
wire i_type_system;
assign i_type_system = opcode == 7'b1110011;
`endif

wire r_type, i_type, s_type, u_type, b_type, j_type;
assign r_type = opcode == 7'b0110011;
`ifdef VIGNA_CORE_ZICSR_EXTENSION
assign i_type = i_type_alu || i_type_jalr || i_type_load || i_type_system;
`else
assign i_type = i_type_alu || i_type_jalr || i_type_load;
`endif
assign s_type = opcode == 7'b0100011;
assign u_type = is_lui || is_auipc;
assign b_type = opcode == 7'b1100011;
assign j_type = opcode == 7'b1101111;

wire [31:0] imm;
assign imm[31]    = effective_inst[31];
assign imm[30:20] = u_type           ? effective_inst[30:20] : {11{effective_inst[31]}};
assign imm[19:12] = u_type || j_type ? effective_inst[19:12] : {8{effective_inst[31]}};
assign imm[11]    = u_type           ? 1'b0 :
                    j_type           ? effective_inst[20] :
                    b_type           ? effective_inst[7] : effective_inst[31];
assign imm[10:5]  = u_type           ? 6'b000000 : effective_inst[30:25];
assign imm[4:1]   = u_type           ? 5'b00000 :
                    u_type           ? 4'b0000 :
                    i_type || j_type ? effective_inst[24:21] : effective_inst[11:8];
assign imm[0]     = i_type           ? effective_inst[20] :
                    s_type           ? effective_inst[7] : 1'b0;


wire [4:0] shamt;
assign shamt = effective_inst[24:20];

//r type
assign is_add  = funct3 == 3'b000 && funct7_zero    && r_type;
assign is_sub  = funct3 == 3'b000 && funct7_sub_sra && r_type;
assign is_sll  = funct3 == 3'b001 && funct7_zero    && r_type;
assign is_slt  = funct3 == 3'b010 && funct7_zero    && r_type;
assign is_sltu = funct3 == 3'b011 && funct7_zero    && r_type;
assign is_xor  = funct3 == 3'b100 && funct7_zero    && r_type;
assign is_srl  = funct3 == 3'b101 && funct7_zero    && r_type;
assign is_sra  = funct3 == 3'b101 && funct7_sub_sra && r_type;
assign is_or   = funct3 == 3'b110 && funct7_zero    && r_type;
assign is_and  = funct3 == 3'b111 && funct7_zero    && r_type;

//i type
assign is_addi  = i_type_alu  && funct3 == 3'b000;
assign is_slli  = i_type_alu  && funct3 == 3'b001;
assign is_slti  = i_type_alu  && funct3 == 3'b010;
assign is_sltiu = i_type_alu  && funct3 == 3'b011;
assign is_xori  = i_type_alu  && funct3 == 3'b100;
assign is_srli  = i_type_alu  && funct3 == 3'b101 && funct7_zero;
assign is_srai  = i_type_alu  && funct3 == 3'b101 && funct7_sub_sra;
assign is_ori   = i_type_alu  && funct3 == 3'b110;
assign is_andi  = i_type_alu  && funct3 == 3'b111;
assign is_jalr  = i_type_jalr && funct3 == 3'b000;
assign is_lb    = i_type_load && funct3 == 3'b000;
assign is_lh    = i_type_load && funct3 == 3'b001;
assign is_lw    = i_type_load && funct3 == 3'b010;
assign is_lbu   = i_type_load && funct3 == 3'b100;
assign is_lhu   = i_type_load && funct3 == 3'b101;

wire is_load;
assign is_load = is_lb || is_lh || is_lw || is_lbu || is_lhu;

//s type
assign is_sb = funct3 == 3'b000 && s_type;
assign is_sh = funct3 == 3'b001 && s_type;
assign is_sw = funct3 == 3'b010 && s_type;

//b type
assign is_beq  = funct3 == 3'b000 && b_type;
assign is_bne  = funct3 == 3'b001 && b_type;
assign is_blt  = funct3 == 3'b100 && b_type;
assign is_bge  = funct3 == 3'b101 && b_type;
assign is_bltu = funct3 == 3'b110 && b_type;
assign is_bgeu = funct3 == 3'b111 && b_type;

//u type
assign is_lui   = opcode == 7'b0110111;
assign is_auipc = opcode == 7'b0010111;

//j type
assign is_jal = j_type;

`ifdef VIGNA_CORE_C_EXTENSION
// C extension instruction decoding
wire [1:0] c_op;
wire [2:0] c_funct3;
wire [4:0] c_rs1, c_rs2, c_rd;
wire [4:0] c_rs1_compressed, c_rs2_compressed; // 3-bit compressed register indices
wire [31:0] c_imm;
wire [31:0] expanded_inst; // Expanded 32-bit instruction from 16-bit C instruction

// Extract C instruction fields
assign c_op = inst[1:0];
assign c_funct3 = inst[15:13];
assign c_rs1 = inst[11:7];
assign c_rs2 = inst[6:2];
assign c_rd = inst[11:7];
assign c_rs1_compressed = {2'b01, inst[9:7]}; // x8-x15 mapping
assign c_rs2_compressed = {2'b01, inst[4:2]}; // x8-x15 mapping

// C instruction type detection
wire c_addi4spn, c_lw, c_sw, c_addi, c_jal, c_li, c_lui, c_srli, c_srai, c_andi, c_sub, c_xor, c_or, c_and;
wire c_j, c_beqz, c_bnez, c_slli, c_lwsp, c_jr, c_mv, c_ebreak, c_jalr, c_add, c_swsp;

// CR format (Compressed Register)
assign c_jr   = (c_op == 2'b10) && (c_funct3 == 3'b100) && (inst[12] == 1'b0) && (inst[6:2] == 5'b00000);
assign c_mv   = (c_op == 2'b10) && (c_funct3 == 3'b100) && (inst[12] == 1'b0) && (inst[6:2] != 5'b00000);
assign c_jalr = (c_op == 2'b10) && (c_funct3 == 3'b100) && (inst[12] == 1'b1) && (inst[6:2] == 5'b00000);
assign c_add  = (c_op == 2'b10) && (c_funct3 == 3'b100) && (inst[12] == 1'b1) && (inst[6:2] != 5'b00000);

// CI format (Compressed Immediate)
assign c_addi = (c_op == 2'b01) && (c_funct3 == 3'b000);
assign c_jal  = (c_op == 2'b01) && (c_funct3 == 3'b001);
assign c_li   = (c_op == 2'b01) && (c_funct3 == 3'b010);
assign c_lui  = (c_op == 2'b01) && (c_funct3 == 3'b011);
assign c_slli = (c_op == 2'b10) && (c_funct3 == 3'b000);
assign c_lwsp = (c_op == 2'b10) && (c_funct3 == 3'b010);

// CSS format (Compressed Stack-relative Store)
assign c_swsp = (c_op == 2'b10) && (c_funct3 == 3'b110);

// CIW format (Compressed Immediate Wide)
assign c_addi4spn = (c_op == 2'b00) && (c_funct3 == 3'b000);

// CL format (Compressed Load)
assign c_lw = (c_op == 2'b00) && (c_funct3 == 3'b010);

// CS format (Compressed Store)
assign c_sw = (c_op == 2'b00) && (c_funct3 == 3'b110);

// CB format (Compressed Branch)
assign c_srli = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b00);
assign c_srai = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b01);
assign c_andi = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b10);
assign c_sub  = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b11) && (inst[6:5] == 2'b00);
assign c_xor  = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b11) && (inst[6:5] == 2'b01);
assign c_or   = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b11) && (inst[6:5] == 2'b10);
assign c_and  = (c_op == 2'b01) && (c_funct3 == 3'b100) && (inst[11:10] == 2'b11) && (inst[6:5] == 2'b11);
assign c_beqz = (c_op == 2'b01) && (c_funct3 == 3'b110);
assign c_bnez = (c_op == 2'b01) && (c_funct3 == 3'b111);

// CJ format (Compressed Jump)
assign c_j = (c_op == 2'b01) && (c_funct3 == 3'b101);

// C instruction immediate generation
wire [31:0] c_imm_addi4spn, c_imm_lw_sw, c_imm_addi, c_imm_jal, c_imm_li, c_imm_lui;
wire [31:0] c_imm_slli, c_imm_lwsp, c_imm_swsp, c_imm_beqz_bnez, c_imm_j;

assign c_imm_addi4spn = {22'b0, inst[10:7], inst[12:11], inst[5], inst[6], 2'b00}; // CIW
assign c_imm_lw_sw = {25'b0, inst[5], inst[12:10], inst[6], 2'b00}; // CL/CS
assign c_imm_addi = {{26{inst[12]}}, inst[12], inst[6:2]}; // CI
assign c_imm_jal = {{20{inst[12]}}, inst[12], inst[8], inst[10:9], inst[6], inst[7], inst[2], inst[11], inst[5:3], 1'b0}; // CJ
assign c_imm_li = {{26{inst[12]}}, inst[12], inst[6:2]}; // CI
assign c_imm_lui = {{14{inst[12]}}, inst[12], inst[6:2], 12'b0}; // CI
assign c_imm_slli = {26'b0, inst[12], inst[6:2]}; // CI
assign c_imm_lwsp = {24'b0, inst[3:2], inst[12], inst[6:4], 2'b00}; // CI
assign c_imm_swsp = {24'b0, inst[8:7], inst[12:9], 2'b00}; // CSS
assign c_imm_beqz_bnez = {{23{inst[12]}}, inst[12], inst[6:5], inst[2], inst[11:10], inst[4:3], 1'b0}; // CB
assign c_imm_j = {{20{inst[12]}}, inst[12], inst[8], inst[10:9], inst[6], inst[7], inst[2], inst[11], inst[5:3], 1'b0}; // CJ

// Expand compressed instructions to 32-bit equivalents
assign expanded_inst = 
    c_addi4spn ? {c_imm_addi4spn[11:0], 5'd2, 3'b000, c_rs2_compressed, 7'b0010011} : // ADDI rd', x2, nzuimm
    c_lw       ? {c_imm_lw_sw[11:0], c_rs1_compressed, 3'b010, c_rs2_compressed, 7'b0000011} : // LW rd', offset(rs1')
    c_sw       ? {c_imm_lw_sw[11:5], c_rs2_compressed, c_rs1_compressed, 3'b010, c_imm_lw_sw[4:0], 7'b0100011} : // SW rs2', offset(rs1')
    c_addi     ? {c_imm_addi[11:0], c_rs1, 3'b000, c_rd, 7'b0010011} : // ADDI rd, rs1, imm
    c_jal      ? {c_imm_jal[20], c_imm_jal[10:1], c_imm_jal[11], c_imm_jal[19:12], 5'd1, 7'b1101111} : // JAL x1, offset
    c_li       ? {c_imm_li[11:0], 5'd0, 3'b000, c_rd, 7'b0010011} : // ADDI rd, x0, imm
    c_lui      ? {c_imm_lui[31:12], c_rd, 7'b0110111} : // LUI rd, imm
    c_srli     ? {7'b0000000, inst[6:2], c_rs1_compressed, 3'b101, c_rs1_compressed, 7'b0010011} : // SRLI rs1', shamt
    c_srai     ? {7'b0100000, inst[6:2], c_rs1_compressed, 3'b101, c_rs1_compressed, 7'b0010011} : // SRAI rs1', shamt
    c_andi     ? {c_imm_addi[11:0], c_rs1_compressed, 3'b111, c_rs1_compressed, 7'b0010011} : // ANDI rs1', imm
    c_sub      ? {7'b0100000, c_rs2_compressed, c_rs1_compressed, 3'b000, c_rs1_compressed, 7'b0110011} : // SUB rs1', rs2'
    c_xor      ? {7'b0000000, c_rs2_compressed, c_rs1_compressed, 3'b100, c_rs1_compressed, 7'b0110011} : // XOR rs1', rs2'
    c_or       ? {7'b0000000, c_rs2_compressed, c_rs1_compressed, 3'b110, c_rs1_compressed, 7'b0110011} : // OR rs1', rs2'
    c_and      ? {7'b0000000, c_rs2_compressed, c_rs1_compressed, 3'b111, c_rs1_compressed, 7'b0110011} : // AND rs1', rs2'
    c_j        ? {c_imm_j[20], c_imm_j[10:1], c_imm_j[11], c_imm_j[19:12], 5'd0, 7'b1101111} : // JAL x0, offset
    c_beqz     ? {c_imm_beqz_bnez[12], c_imm_beqz_bnez[10:5], 5'd0, c_rs1_compressed, 3'b000, c_imm_beqz_bnez[4:1], c_imm_beqz_bnez[11], 7'b1100011} : // BEQ rs1', x0, offset
    c_bnez     ? {c_imm_beqz_bnez[12], c_imm_beqz_bnez[10:5], 5'd0, c_rs1_compressed, 3'b001, c_imm_beqz_bnez[4:1], c_imm_beqz_bnez[11], 7'b1100011} : // BNE rs1', x0, offset
    c_slli     ? {7'b0000000, inst[6:2], c_rs1, 3'b001, c_rd, 7'b0010011} : // SLLI rd, rs1, shamt
    c_lwsp     ? {c_imm_lwsp[11:0], 5'd2, 3'b010, c_rd, 7'b0000011} : // LW rd, offset(x2)
    c_jr       ? {12'b0, c_rs1, 3'b000, 5'd0, 7'b1100111} : // JALR x0, 0(rs1)
    c_mv       ? {7'b0000000, c_rs2, 5'd0, 3'b000, c_rd, 7'b0110011} : // ADD rd, x0, rs2
    c_jalr     ? {12'b0, c_rs1, 3'b000, 5'd1, 7'b1100111} : // JALR x1, 0(rs1)
    c_add      ? {7'b0000000, c_rs2, c_rs1, 3'b000, c_rd, 7'b0110011} : // ADD rd, rs1, rs2
    c_swsp     ? {c_imm_swsp[11:5], c_rs2, 5'd2, 3'b010, c_imm_swsp[4:0], 7'b0100011} : // SW rs2, offset(x2)
    32'h00000013; // Default to NOP (ADDI x0, x0, 0)

// Select between original 32-bit instruction and expanded C instruction
wire [31:0] effective_inst;
assign effective_inst = (inst_is_16bit) ? expanded_inst : inst;
`else
wire [31:0] effective_inst;
assign effective_inst = inst;
`endif

`ifdef VIGNA_CORE_M_EXTENSION
//m type
wire is_m_coproc;
assign is_m_coproc = r_type && funct7 == 7'b0000001;
`endif

`ifdef VIGNA_CORE_ZICSR_EXTENSION
//csr type (system instructions)
wire is_csrrw, is_csrrs, is_csrrc, is_csrrwi, is_csrrsi, is_csrrci;
assign is_csrrw  = i_type_system && funct3 == 3'b001;
assign is_csrrs  = i_type_system && funct3 == 3'b010;
assign is_csrrc  = i_type_system && funct3 == 3'b011;
assign is_csrrwi = i_type_system && funct3 == 3'b101;
assign is_csrrsi = i_type_system && funct3 == 3'b110;
assign is_csrrci = i_type_system && funct3 == 3'b111;

`ifdef VIGNA_CORE_INTERRUPT
// MRET instruction (Machine Return from trap)
wire is_mret;
assign is_mret = i_type_system && funct3 == 3'b000 && rs2 == 5'b00010 && rd == 5'b00000 && rs1 == 5'b00000;
`endif

wire is_csr_op;
assign is_csr_op = is_csrrw || is_csrrs || is_csrrc || is_csrrwi || is_csrrsi || is_csrrci
`ifdef VIGNA_CORE_INTERRUPT
                   || is_mret
`endif
                   ;
`endif

//rs1 from reg
wire [31:0] rs1_val;
//rs2 from reg
wire [31:0] rs2_val;

//cpu regs
`ifdef VIGNA_CORE_E_EXTENSION
    reg [31:0] cpu_regs[15:1];
    assign rs1_val = rs1 == 0 ? 32'd0 : cpu_regs[rs1[3:0]];
    assign rs2_val = rs2 == 0 ? 32'd0 : cpu_regs[rs2[3:0]];
`else
    reg [31:0] cpu_regs[31:1];
    assign rs1_val = rs1 == 0 ? 32'd0 : cpu_regs[rs1];
    assign rs2_val = rs2 == 0 ? 32'd0 : cpu_regs[rs2];
`endif

`ifdef VIGNA_CORE_ZICSR_EXTENSION
//csr regs - implementing basic set for now
reg [31:0] csr_regs[4095:0];  // Full CSR address space
wire [11:0] csr_addr;
assign csr_addr = imm[11:0];  // CSR address is in immediate field

// CSR read value
wire [31:0] csr_rval;
assign csr_rval = csr_regs[csr_addr];

`ifdef VIGNA_CORE_INTERRUPT
// Machine-level interrupt CSR addresses (RISC-V standard)
localparam [11:0] CSR_MSTATUS  = 12'h300;  // Machine status
localparam [11:0] CSR_MIE      = 12'h304;  // Machine interrupt enable
localparam [11:0] CSR_MTVEC    = 12'h305;  // Machine trap vector base address
localparam [11:0] CSR_MSCRATCH = 12'h340;  // Machine scratch register
localparam [11:0] CSR_MEPC     = 12'h341;  // Machine exception program counter
localparam [11:0] CSR_MCAUSE   = 12'h342;  // Machine cause register
localparam [11:0] CSR_MTVAL    = 12'h343;  // Machine trap value
localparam [11:0] CSR_MIP      = 12'h344;  // Machine interrupt pending

// Interrupt control signals
reg interrupt_taken;
reg [31:0] interrupt_cause;
wire [31:0] mstatus, mie, mip, mtvec, mepc, mcause, mtval, mscratch;
assign mstatus  = csr_regs[CSR_MSTATUS];
assign mie      = csr_regs[CSR_MIE];
assign mip      = csr_regs[CSR_MIP];
assign mtvec    = csr_regs[CSR_MTVEC];
assign mepc     = csr_regs[CSR_MEPC];
assign mcause   = csr_regs[CSR_MCAUSE];
assign mtval    = csr_regs[CSR_MTVAL];
assign mscratch = csr_regs[CSR_MSCRATCH];

// Interrupt pending bits (updated by hardware)
wire [2:0] irq_pending;
assign irq_pending = {ext_irq, timer_irq, soft_irq};

// Global interrupt enable from mstatus.MIE (bit 3)
wire global_irq_enable;
assign global_irq_enable = mstatus[3];

// Check for pending and enabled interrupts
wire ext_irq_ready, timer_irq_ready, soft_irq_ready;
assign ext_irq_ready   = irq_pending[2] & mie[11] & global_irq_enable; // MEI
assign timer_irq_ready = irq_pending[1] & mie[7]  & global_irq_enable; // MTI  
assign soft_irq_ready  = irq_pending[0] & mie[3]  & global_irq_enable; // MSI

// Interrupt request (prioritized: external > timer > software)
wire interrupt_request;
assign interrupt_request = ext_irq_ready | timer_irq_ready | soft_irq_ready;
`endif
`endif

wire [31:0] op1, op2;
`ifdef VIGNA_CORE_ZICSR_EXTENSION
assign op1 = is_jal || u_type   ? imm : 
             is_csr_op          ? csr_rval : rs1_val;
assign op2 = (r_type || b_type)   ? rs2_val :
             (is_auipc || j_type) ? inst_addr :
             (is_slli || is_srli) ? {27'b0, shamt} :
             is_lui               ? 32'd0 :
             is_csr_op            ? ((is_csrrwi || is_csrrsi || is_csrrci) ? {27'b0, rs1} : rs1_val) :
             imm;
`else
assign op1 = is_jal || u_type   ? imm : rs1_val;
assign op2 = (r_type || b_type)   ? rs2_val :
             (is_auipc || j_type) ? inst_addr :
             (is_slli || is_srli) ? {27'b0, shamt} :
             is_lui               ? 32'd0 : imm; 
`endif 

//backend state
reg [3:0] exec_state;

//source regex_jump
reg [31:0] d1, d2, d3;

//result
wire [31:0] dr;

//write back
`ifdef VIGNA_CORE_E_EXTENSION
    reg [3:0] wb_reg;
`else
    reg [4:0] wb_reg;
`endif 

    reg [4:0] shift_cnt;
    reg [2:0] l_sll_srl_sra;
    wire [31:0] shift_val;
    wire is_shift;
    assign is_shift = is_sll || is_slli || is_srl || is_srli || is_sra || is_srai;
`ifdef VIGNA_CORE_TWO_STAGE_SHIFT
    wire first_shift_stage;
    assign first_shift_stage = shift_cnt[4:2] != 0;
`endif

wire cmp_eq;
wire abs_lt;
wire signed_lt;
wire unsigned_lt;
assign cmp_eq      = d1 == d2;
assign abs_lt      = d1[30:0] < d2[30:0];
assign signed_lt   = (d1[31] ^ d2[31]) ? d1[31] : abs_lt;
assign unsigned_lt = (d1[31] ^ d2[31]) ? d2[31] : abs_lt;

wire [31:0] add_result;
`ifdef VIGNA_CORE_PRELOAD_NEGATIVE
assign add_result = d1 + d2 + is_sub;
`else
assign add_result = d1 + (is_sub ? {~d2 + 32'd1} : d2);
`endif

//alu comb logic
assign dr = 
    is_add || is_addi || is_jal || s_type
     || is_jalr || is_load || u_type
     || is_sub                      ? add_result : 
    is_slt || is_slti || is_blt     ? {31'd0, signed_lt} :
    is_bge                          ? {31'd0, ~signed_lt} :
    is_sltu || is_sltiu || is_bltu  ? {31'd0, unsigned_lt} : 
    is_bgeu                         ? {31'd0, ~unsigned_lt} :
    is_xor || is_xori               ? d1 ^ d2 :  
    is_or || is_ori                 ? d1 | d2 : 
    is_and || is_andi               ? d1 & d2 : 
    is_beq                          ? {31'd0, cmp_eq} : 
    is_bne                          ? {31'd0, ~cmp_eq} : 32'd0;

assign shift_val =
`ifdef  VIGNA_CORE_TWO_STAGE_SHIFT
    l_sll_srl_sra[2]  ? (first_shift_stage ? {d3[27:0], 4'b0000} : {d3[30:0], 1'b0}) :
    l_sll_srl_sra[1]  ? (first_shift_stage ? {4'b0000, d3[31:4]} : {1'b0, d3[31:1]}) :
    l_sll_srl_sra[0]  ? (first_shift_stage ? {{4{d3[31]}}, d3[31:4]} : {d3[31], d3[31:1]}) : 32'd0;
`else 
    l_sll_srl_sra[2]  ? {d3[30:0], 1'b0} :
    l_sll_srl_sra[1]  ? {1'b0, d3[31:1]} :
    l_sll_srl_sra[0]  ? {d3[31], d3[31:1]} : 32'd0;
`endif

wire [31:0] inst_add_result;
`ifdef VIGNA_CORE_C_EXTENSION
wire [31:0] pc_increment;
assign pc_increment = inst_is_16bit ? 32'd2 : 32'd4;
assign inst_add_result = inst_addr + (b_type ? imm : pc_increment);
`else
assign inst_add_result = inst_addr + (b_type ? imm : 32'd4);
`endif

reg ex_branch;
reg ex_jump;
reg [3:0] ex_type;
reg [3:0] ls_strb;
reg ls_sign_extend;

assign pc_next =  interrupt_taken     ? interrupt_cause :
                  `ifdef VIGNA_CORE_INTERRUPT
                  (ex_jump && is_mret)  ? mepc :
                  `endif
                  ex_jump           ? dr :
                  ex_branch & dr[0] ? d3 : 
                  `ifdef VIGNA_CORE_C_EXTENSION
                  pc + pc_increment;
                  `else
                  pc + 32'd4;
                  `endif

reg write_mem;

wire is_jump = is_jal || is_jalr;

`ifdef VIGNA_CORE_M_EXTENSION
    reg m_valid;
    wire m_ready;
    wire [31:0] m_result;
    vigna_m_ext mul_unit(
        .clk(clk),
        .resetn(resetn),
        .valid(m_valid),
        .ready(m_ready),
        .op1(d1),
        .op2(d2),
        .result(m_result),
        .func(d3[2:0])
    );
`endif


//part2. executon unit
always @ (posedge clk) begin
    //reset logic
    if (!resetn) begin
        d_valid        <= 0;
        d_addr         <= 0;
        d_wdata        <= 0;
        d_wstrb        <= 0;
        d1             <= 0;
        d2             <= 0;
        d3             <= 0;
        exec_state     <= 0;
        wb_reg         <= 0;
        ex_jump        <= 0;
        `ifdef VIGNA_CORE_ZICSR_EXTENSION
        // Initialize CSR registers to 0  
        for (integer i = 0; i < 4096; i = i + 1) begin
            csr_regs[i] <= 32'h00000000;
        end
        `ifdef VIGNA_CORE_INTERRUPT
        // Initialize interrupt-specific CSRs with minimal changes
        // Keep mstatus at 0 for compatibility with existing tests
        csr_regs[CSR_MIE]     <= 32'h00000000; // All interrupts disabled
        csr_regs[CSR_MIP]     <= 32'h00000000; // No pending interrupts
        csr_regs[CSR_MTVEC]   <= 32'h00000000; // Trap vector at address 0
        `endif
        `endif
        ex_branch      <= 0;
        write_mem      <= 0;
        ls_strb        <= 0;
        ls_sign_extend <= 0;
        // Reset all CPU registers to 0
        `ifdef VIGNA_CORE_E_EXTENSION
            for (integer i = 1; i <= 15; i = i + 1)
                cpu_regs[i] <= 32'd0;
        `else
            for (integer i = 1; i <= 31; i = i + 1)
                cpu_regs[i] <= 32'd0;
        `endif
        
        `ifdef VIGNA_CORE_STACK_ADDR_RESET_ENABLE
            cpu_regs[2] <= `VIGNA_CORE_STACK_ADDR_RESET_VALUE;
        `endif
        shift_cnt <= 0;
        l_sll_srl_sra <= 0;
        `ifdef VIGNA_CORE_INTERRUPT
        interrupt_taken <= 0;
        interrupt_cause <= 0;
        `endif
    end else begin
        `ifdef VIGNA_CORE_INTERRUPT
        // Update interrupt pending register based on external signals
        csr_regs[CSR_MIP][11] <= ext_irq;    // MEI - Machine External Interrupt
        csr_regs[CSR_MIP][7]  <= timer_irq;  // MTI - Machine Timer Interrupt  
        csr_regs[CSR_MIP][3]  <= soft_irq;   // MSI - Machine Software Interrupt
        
        // Check for interrupt request during instruction fetch
        if (exec_state == 4'b0000 && fetched && interrupt_request && !interrupt_taken) begin
            // Take interrupt: save state and jump to handler
            interrupt_taken <= 1;
            csr_regs[CSR_MEPC] <= pc; // Save current PC
            csr_regs[CSR_MSTATUS][7] <= mstatus[3]; // Save current MIE to MPIE
            csr_regs[CSR_MSTATUS][3] <= 0; // Disable interrupts (clear MIE)
            
            // Determine interrupt cause and set mcause
            if (ext_irq_ready) begin
                csr_regs[CSR_MCAUSE] <= 32'h80000000 | 32'd11; // External interrupt
                interrupt_cause <= mtvec; // Jump to trap handler
            end else if (timer_irq_ready) begin
                csr_regs[CSR_MCAUSE] <= 32'h80000000 | 32'd7;  // Timer interrupt
                interrupt_cause <= mtvec; // Jump to trap handler
            end else if (soft_irq_ready) begin
                csr_regs[CSR_MCAUSE] <= 32'h80000000 | 32'd3;  // Software interrupt
                interrupt_cause <= mtvec; // Jump to trap handler
            end
        end else begin
            interrupt_taken <= 0;
        end
        `endif
        
        //state machine
        case (exec_state)
            4'b0000: begin
                if (fetched) begin
                    d1 <= op1;
                    `ifdef VIGNA_CORE_PRELOAD_NEGATIVE
                    d2 <= (is_sub ? ~op2 : op2);
                    `else
                    d2 <= op2;
                    `endif
                    if (s_type) begin
                        d3 <= rs2_val;
                    end else if (b_type) begin
                        d3 <= inst_add_result;
                    end else if (is_jal || is_jalr) begin
                        d3 <= inst_add_result;
                    end else if (is_shift) begin
                        l_sll_srl_sra <= {is_sll || is_slli, is_srl || is_srli, is_sra || is_srai};
                        d3 <= op1;
                        shift_cnt <= op2[4:0];
                    `ifdef VIGNA_CORE_M_EXTENSION
                    end else if (is_m_coproc) begin 
                        d3[2:0] <= funct3;
                        m_valid   <= 1;
                    `endif
                    end
                                    
                    if (u_type || j_type || i_type || r_type) begin
                        `ifdef VIGNA_CORE_E_EXTENSION
                            wb_reg <= rd[3:0];
                        `else 
                            wb_reg <= rd;
                        `endif
                    end else begin
                        wb_reg <= 0;
                    end
                    ex_branch   <= b_type;
                    ex_jump     <= is_jal || is_jalr;

                    //next state logic
                    if (is_load || s_type) begin
                        exec_state <= 4'b0001;
                        write_mem <= is_load ? 1'b0 : 1'b1;
                    end
                    else if (is_jal || is_jalr) begin
                        exec_state <= 4'b0100;
                    end
                    else if (b_type) begin
                        exec_state <= 4'b1000;
                    end
                    else if (is_shift) begin
                        exec_state <= 4'b0110;
                    end
                    `ifdef VIGNA_CORE_M_EXTENSION
                    else if (is_m_coproc) begin
                        exec_state <= 4'b1001;
                    end
                    `endif
                    `ifdef VIGNA_CORE_ZICSR_EXTENSION
                    else if (is_csr_op) begin
                        exec_state <= 4'b1010;
                    end
                    `endif 
                    else begin
                        exec_state <= 4'b0010;
                    end

                    //set strobe
                    if (is_lw || is_sw) ls_strb <= 4'b1111;
                    else if (is_lh || is_lhu || is_sh) ls_strb <= 4'b0011;
                    else if (is_lb || is_lbu || is_sb) ls_strb <= 4'b0001;

                    if (is_lw || is_lh || is_lb) ls_sign_extend <= 1;
                    else ls_sign_extend <= 0;
                end
            end
            4'b0001: begin
                //load/store func
                if (!write_mem) begin
                    d_valid    <= 1;
                    `ifdef VIGNA_CORE_ALIGNMENT 
                        d_addr <= dr & 32'hfffffffc;
                        shift_cnt <= dr[1:0];
                    `else
                        d_addr <= dr;  
                    `endif
                    d_wstrb    <= 0;
                    exec_state <= 4'b0011;
                end else begin
                    d_valid    <= 1;
                    `ifdef VIGNA_CORE_ALIGNMENT 
                        d_addr <= dr & 32'hfffffffc;
                        shift_cnt[1:0] <= dr[1:0];
                        d_wdata    <= d3 << ({3'b000, dr[1:0]} << 3);
                        d_wstrb    <= ls_strb << dr[1:0];
                    `else
                        d_addr <= dr;  
                        d_wdata    <= d3;
                        d_wstrb    <= ls_strb;
                    `endif
                    exec_state <= 4'b0101;
                end
            end
            4'b0010: begin
                //calc func
                exec_state <= 0;
                if (wb_reg != 0) begin
                    cpu_regs[wb_reg] <= dr;
                end
            end
            4'b0100: begin
                //jump func
                exec_state <= 0;
                ex_jump    <= 0;
                if (wb_reg != 0) begin
                    cpu_regs[wb_reg] <= d3;
                end
            end
            4'b1000: begin
                //branch func
                exec_state     <= 0;
                ex_branch      <= 0;
            end
            4'b0011: begin
                //load wait stage
                if (d_ready) begin
                    exec_state <= 0;
                    d_valid    <= 0;
                    if (wb_reg != 0) begin
                        `ifdef VIGNA_CORE_ALIGNMENT
                            case ({shift_cnt[1:0], ls_strb})
                                6'b000001: cpu_regs[wb_reg] <= {ls_sign_extend ? {24{d_rdata[ 7]}} : 24'd0, d_rdata[ 7: 0]};
                                6'b010001: cpu_regs[wb_reg] <= {ls_sign_extend ? {24{d_rdata[15]}} : 24'd0, d_rdata[15: 8]};
                                6'b100001: cpu_regs[wb_reg] <= {ls_sign_extend ? {24{d_rdata[23]}} : 24'd0, d_rdata[23:16]};
                                6'b110001: cpu_regs[wb_reg] <= {ls_sign_extend ? {24{d_rdata[31]}} : 24'd0, d_rdata[31:24]};
                                6'b000011: cpu_regs[wb_reg] <= {ls_sign_extend ? {16{d_rdata[15]}} : 16'd0, d_rdata[15: 0]};
                                6'b100011: cpu_regs[wb_reg] <= {ls_sign_extend ? {16{d_rdata[31]}} : 16'd0, d_rdata[31:16]};
                                6'b001111: cpu_regs[wb_reg] <= d_rdata;
                                default: cpu_regs[wb_reg] <= 32'd0;
                            endcase
                        `else 
                            if      (!ls_sign_extend)    cpu_regs[wb_reg] <= d_rdata & {{8{ls_strb[3]}}, {8{ls_strb[2]}}, {8{ls_strb[1]}}, {8{ls_strb[0]}}};
                            else if (ls_strb == 4'b0001) cpu_regs[wb_reg] <= {{24{d_rdata[7]}}, d_rdata[7:0]};
                            else if (ls_strb == 4'b0011) cpu_regs[wb_reg] <= {{16{d_rdata[15]}}, d_rdata[15:0]};
                            else                         cpu_regs[wb_reg] <= d_rdata;
                        `endif      
                    end
                end
            end
            4'b0101: begin
                //store wait stage
                if (d_ready) begin
                    exec_state <= 0;
                    d_valid    <= 0;
                    d_wstrb    <= 4'd0;
                    d_wdata    <= 0;
                end
            end
            4'b0110: begin
                //shift func
                if (shift_cnt == 0) begin
                    exec_state <= 0;
                    cpu_regs[wb_reg] <= d3;
                end else begin
                    `ifdef VIGNA_CORE_TWO_STAGE_SHIFT
                    if (first_shift_stage)
                        shift_cnt <= shift_cnt - 4;
                    else
                    `endif
                        shift_cnt <= shift_cnt - 1;
                    d3 <= shift_val;
                end
            end 
            `ifdef VIGNA_CORE_M_EXTENSION
            4'b1001: begin
                m_valid <= 0;
                if (m_ready) begin
                    cpu_regs[wb_reg] <= m_result;
                    exec_state <= 0;
                end
            end
            `endif
            `ifdef VIGNA_CORE_ZICSR_EXTENSION
            4'b1010: begin
                //csr operation
                exec_state <= 0;
                `ifdef VIGNA_CORE_INTERRUPT
                if (is_mret) begin
                    // Machine return: restore PC and interrupt enable
                    // This will be handled in pc_next logic
                    csr_regs[CSR_MSTATUS][3] <= mstatus[7]; // Restore MIE from MPIE
                    csr_regs[CSR_MSTATUS][7] <= 1; // Set MPIE to 1
                    ex_jump <= 1; // Jump to MEPC
                end else begin
                `endif
                    if (wb_reg != 0) begin
                        cpu_regs[wb_reg] <= op1;  // write old CSR value to rd
                    end
                    // Update CSR based on operation type
                    if (is_csrrw || is_csrrwi) begin
                        // CSR = rs1_val or imm
                        csr_regs[csr_addr] <= op2;
                    end
                    else if (is_csrrs || is_csrrsi) begin
                        // CSR = CSR | (rs1_val or imm)
                        if (rs1 != 0) begin // only write if rs1 != 0
                            csr_regs[csr_addr] <= op1 | op2;
                        end
                    end
                    else if (is_csrrc || is_csrrci) begin
                        // CSR = CSR & ~(rs1_val or imm)
                        if (rs1 != 0) begin // only write if rs1 != 0
                            csr_regs[csr_addr] <= op1 & ~op2;
                        end
                    end
                `ifdef VIGNA_CORE_INTERRUPT
                end
                `endif
            end
            `endif
            default: begin
                exec_state <= 0;
            end
        endcase
    end
end

wire is_branch;
assign is_branch = is_beq || is_bne || is_blt || is_bge || is_bltu || is_bgeu;

assign fetch_received = (exec_state == 4'b0000 && !is_jump && !is_branch)
                        || (exec_state == 4'b0100)
                        || (exec_state == 4'b1000)
                        `ifdef VIGNA_CORE_ZICSR_EXTENSION
                        || (exec_state == 4'b1010)
                        `endif
                        ;

endmodule

`endif
